// Implement module called full_adder