module light(
    // Declare downstairs and upstairs input
    // Declare stair light output
);

    // Enter logic equation here

endmodule